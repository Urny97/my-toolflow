-- David Leifker    
-- 128bit AES Encryption Implementation
-- Contains code for sbox tables lookup for subbytes function
-- Filename: bytesub.vhd

library ieee;
use ieee.std_logic_1164.all;

entity AES_sbox is
  port( SB_in :in std_logic_vector( 7 downto 0 );
    SB_out :out std_logic_vector( 7 downto 0 )
  );
end AES_sbox;

architecture Behavioral of AES_sbox is

begin
  process(SB_in)
  begin
    case SB_in is
    when "01000010" => SB_out <=  "00101100";
    when "10101000" => SB_out <=  "11000010";
    when "10110110" => SB_out <=  "01001110";
    when "00011010" => SB_out <=  "10100010";
    when "00111000" => SB_out <=  "00000111";
    when "11011000" => SB_out <=  "01100001";
    when "00000101" => SB_out <=  "01101011";
    when "00101111" => SB_out <=  "00010101";
    when "00110101" => SB_out <=  "10010110";
    when "00111111" => SB_out <=  "01110101";
    when "10000010" => SB_out <=  "00010011";
    when "00000110" => SB_out <=  "01101111";
    when "00100011" => SB_out <=  "00100110";
    when "10010010" => SB_out <=  "01001111";
    when "11000000" => SB_out <=  "10111010";
    when "11010000" => SB_out <=  "01110000";
    when "10111010" => SB_out <=  "11110100";
    when "10010111" => SB_out <=  "10001000";
    when "10101011" => SB_out <=  "01100010";
    when "11100110" => SB_out <=  "10001110";
    when "11101100" => SB_out <=  "11001110";
    when "00011101" => SB_out <=  "10100100";
    when "00000000" => SB_out <=  "01100011";
    when "10100010" => SB_out <=  "00111010";
    when "11000001" => SB_out <=  "01111000";
    when "00011001" => SB_out <=  "11010100";
    when "01101110" => SB_out <=  "10011111";
    when "11101011" => SB_out <=  "11101001";
    when "11101111" => SB_out <=  "11011111";
    when "00100111" => SB_out <=  "11001100";
    when "11110100" => SB_out <=  "10111111";
    when "00000001" => SB_out <=  "01111100";
    when "00011011" => SB_out <=  "10101111";
    when "01110111" => SB_out <=  "11110101";
    when "11010101" => SB_out <=  "00000011";
    when "00010111" => SB_out <=  "11110000";
    when "00111100" => SB_out <=  "11101011";
    when "10111011" => SB_out <=  "11101010";
    when "01000000" => SB_out <=  "00001001";
    when "11111011" => SB_out <=  "00001111";
    when "01111001" => SB_out <=  "10110110";
    when "10110000" => SB_out <=  "11100111";
    when "10100100" => SB_out <=  "01001001";
    when "11000010" => SB_out <=  "00100101";
    when "11110111" => SB_out <=  "01101000";
    when "00110100" => SB_out <=  "00011000";
    when "01011100" => SB_out <=  "01001010";
    when "00001101" => SB_out <=  "11010111";
    when "00111110" => SB_out <=  "10110010";
    when "01010010" => SB_out <=  "00000000";
    when "01001111" => SB_out <=  "10000100";
    when "11000101" => SB_out <=  "10100110";
    when "11110110" => SB_out <=  "01000010";
    when "01110110" => SB_out <=  "00111000";
    when "00100010" => SB_out <=  "10010011";
    when "00101011" => SB_out <=  "11110001";
    when "11001000" => SB_out <=  "11101000";
    when "01010110" => SB_out <=  "10110001";
    when "10101111" => SB_out <=  "01111001";
    when "11011010" => SB_out <=  "01010111";
    when "11111010" => SB_out <=  "00101101";
    when "00101110" => SB_out <=  "00110001";
    when "11011001" => SB_out <=  "00110101";
    when "11100000" => SB_out <=  "11100001";
    when "01101111" => SB_out <=  "10101000";
    when "11100100" => SB_out <=  "01101001";
    when "01000101" => SB_out <=  "01101110";
    when "00001000" => SB_out <=  "00110000";
    when "00000010" => SB_out <=  "01110111";
    when "00011000" => SB_out <=  "10101101";
    when "00010100" => SB_out <=  "11111010";
    when "01000001" => SB_out <=  "10000011";
    when "10101110" => SB_out <=  "11100100";
    when "10100110" => SB_out <=  "00100100";
    when "01110000" => SB_out <=  "01010001";
    when "01010100" => SB_out <=  "00100000";
    when "11100001" => SB_out <=  "11111000";
    when "10111000" => SB_out <=  "01101100";
    when "00100110" => SB_out <=  "11110111";
    when "10110011" => SB_out <=  "01101101";
    when "11000100" => SB_out <=  "00011100";
    when "11100111" => SB_out <=  "10010100";
    when "11101010" => SB_out <=  "10000111";
    when "00001100" => SB_out <=  "11111110";
    when "00110110" => SB_out <=  "00000101";
    when "01010000" => SB_out <=  "01010011";
    when "11101000" => SB_out <=  "10011011";
    when "10001110" => SB_out <=  "00011001";
    when "11001001" => SB_out <=  "11011101";
    when "11001011" => SB_out <=  "00011111";
    when "10111100" => SB_out <=  "01100101";
    when "00100100" => SB_out <=  "00110110";
    when "01011110" => SB_out <=  "01011000";
    when "01001000" => SB_out <=  "01010010";
    when "10000011" => SB_out <=  "11101100";
    when "11100101" => SB_out <=  "11011001";
    when "11011101" => SB_out <=  "11000001";
    when "00010000" => SB_out <=  "11001010";
    when "01001101" => SB_out <=  "11100011";
    when "01111010" => SB_out <=  "11011010";
    when "11010100" => SB_out <=  "01001000";
    when "00101100" => SB_out <=  "01110001";
    when "01011011" => SB_out <=  "00111001";
    when "01011101" => SB_out <=  "01001100";
    when "10011100" => SB_out <=  "11011110";
    when "01001110" => SB_out <=  "00101111";
    when "11001110" => SB_out <=  "10001011";
    when "00011111" => SB_out <=  "11000000";
    when "00101010" => SB_out <=  "11100101";
    when "11110000" => SB_out <=  "10001100";
    when "00110111" => SB_out <=  "10011010";
    when "11101101" => SB_out <=  "01010101";
    when "11100011" => SB_out <=  "00010001";
    when "10011011" => SB_out <=  "00010100";
    when "01010001" => SB_out <=  "11010001";
    when "10100101" => SB_out <=  "00000110";
    when "01011111" => SB_out <=  "11001111";
    when "01100001" => SB_out <=  "11101111";
    when "10001010" => SB_out <=  "01111110";
    when "00101001" => SB_out <=  "10100101";
    when "00110000" => SB_out <=  "00000100";
    when "01100111" => SB_out <=  "10000101";
    when "10101100" => SB_out <=  "10010001";
    when "11010010" => SB_out <=  "10110101";
    when "00100000" => SB_out <=  "10110111";
    when "10000101" => SB_out <=  "10010111";
    when "01101001" => SB_out <=  "11111001";
    when "00000100" => SB_out <=  "11110010";
    when "10110100" => SB_out <=  "10001101";
    when "01100010" => SB_out <=  "10101010";
    when "01101010" => SB_out <=  "00000010";
    when "01000111" => SB_out <=  "10100000";
    when "00111001" => SB_out <=  "00010010";
    when "11010001" => SB_out <=  "00111110";
    when "10010011" => SB_out <=  "11011100";
    when "10011101" => SB_out <=  "01011110";
    when "01110101" => SB_out <=  "10011101";
    when "11001111" => SB_out <=  "10001010";
    when "00001011" => SB_out <=  "00101011";
    when "01111111" => SB_out <=  "11010010";
    when "11010011" => SB_out <=  "01100110";
    when "00011100" => SB_out <=  "10011100";
    when "11111110" => SB_out <=  "10111011";
    when "00011110" => SB_out <=  "01110010";
    when "10000001" => SB_out <=  "00001100";
    when "10001011" => SB_out <=  "00111101";
    when "00010110" => SB_out <=  "01000111";
    when "10010100" => SB_out <=  "00100010";
    when "10110101" => SB_out <=  "11010101";
    when "01110011" => SB_out <=  "10001111";
    when "11011111" => SB_out <=  "10011110";
    when "11111001" => SB_out <=  "10011001";
    when "10101010" => SB_out <=  "10101100";
    when "10111101" => SB_out <=  "01111010";
    when "11000111" => SB_out <=  "11000110";
    when "11110010" => SB_out <=  "10001001";
    when "01101000" => SB_out <=  "01000101";
    when "10010000" => SB_out <=  "01100000";
    when "00110001" => SB_out <=  "11000111";
    when "01011000" => SB_out <=  "01101010";
    when "10000000" => SB_out <=  "11001101";
    when "10000100" => SB_out <=  "01011111";
    when "10001111" => SB_out <=  "01110011";
    when "10110111" => SB_out <=  "10101001";
    when "10011000" => SB_out <=  "01000110";
    when "01111101" => SB_out <=  "11111111";
    when "10000111" => SB_out <=  "00010111";
    when "11110101" => SB_out <=  "11100110";
    when "11000110" => SB_out <=  "10110100";
    when "10110010" => SB_out <=  "00110111";
    when "01101011" => SB_out <=  "01111111";
    when "01111100" => SB_out <=  "00010000";
    when "10110001" => SB_out <=  "11001000";
    when "00111011" => SB_out <=  "11100010";
    when "01000100" => SB_out <=  "00011011";
    when "11111111" => SB_out <=  "00010110";
    when "01100110" => SB_out <=  "00110011";
    when "01111110" => SB_out <=  "11110011";
    when "10100001" => SB_out <=  "00110010";
    when "00101101" => SB_out <=  "11011000";
    when "01011010" => SB_out <=  "10111110";
    when "00111101" => SB_out <=  "00100111";
    when "10101101" => SB_out <=  "10010101";
    when "10000110" => SB_out <=  "01000100";
    when "00010010" => SB_out <=  "11001001";
    when "11110001" => SB_out <=  "10100001";
    when "01101101" => SB_out <=  "00111100";
    when "10011010" => SB_out <=  "10111000";
    when "01000110" => SB_out <=  "01011010";
    when "01001001" => SB_out <=  "00111011";
    when "10100000" => SB_out <=  "11100000";
    when "11101110" => SB_out <=  "00101000";
    when "11111101" => SB_out <=  "01010100";
    when "00001111" => SB_out <=  "01110110";
    when "00111010" => SB_out <=  "10000000";
    when "11100010" => SB_out <=  "10011000";
    when "01110001" => SB_out <=  "10100011";
    when "11111000" => SB_out <=  "01000001";
    when "11000011" => SB_out <=  "00101110";
    when "00010101" => SB_out <=  "01011001";
    when "01010011" => SB_out <=  "11101101";
    when "01110010" => SB_out <=  "01000000";
    when "10111110" => SB_out <=  "10101110";
    when "00001110" => SB_out <=  "10101011";
    when "00010001" => SB_out <=  "10000010";
    when "10001100" => SB_out <=  "01100100";
    when "01001010" => SB_out <=  "11010110";
    when "10101001" => SB_out <=  "11010011";
    when "11001100" => SB_out <=  "01001011";
    when "10001101" => SB_out <=  "01011101";
    when "11001010" => SB_out <=  "01110100";
    when "10001001" => SB_out <=  "10100111";
    when "10010001" => SB_out <=  "10000001";
    when "11011011" => SB_out <=  "10111001";
    when "00010011" => SB_out <=  "01111101";
    when "00100101" => SB_out <=  "00111111";
    when "01100000" => SB_out <=  "11010000";
    when "01001100" => SB_out <=  "00101001";
    when "10011111" => SB_out <=  "11011011";
    when "11101001" => SB_out <=  "00011110";
    when "00001001" => SB_out <=  "00000001";
    when "00000111" => SB_out <=  "11000101";
    when "01011001" => SB_out <=  "11001011";
    when "01111011" => SB_out <=  "00100001";
    when "10001000" => SB_out <=  "11000100";
    when "10111111" => SB_out <=  "00001000";
    when "00101000" => SB_out <=  "00110100";
    when "10100111" => SB_out <=  "01011100";
    when "10111001" => SB_out <=  "01010110";
    when "00000011" => SB_out <=  "01111011";
    when "00110010" => SB_out <=  "00100011";
    when "01001011" => SB_out <=  "10110011";
    when "11110011" => SB_out <=  "00001101";
    when "01010111" => SB_out <=  "01011011";
    when "11011100" => SB_out <=  "10000110";
    when "10010101" => SB_out <=  "00101010";
    when "10010110" => SB_out <=  "10010000";
    when "01100011" => SB_out <=  "11111011";
    when "01100101" => SB_out <=  "01001101";
    when "11010111" => SB_out <=  "00001110";
    when "01110100" => SB_out <=  "10010010";
    when "11001101" => SB_out <=  "10111101";
    when "01010101" => SB_out <=  "11111100";
    when "01101100" => SB_out <=  "01010000";
    when "10100011" => SB_out <=  "00001010";
    when "11111100" => SB_out <=  "10110000";
    when "10011110" => SB_out <=  "00001011";
    when "11011110" => SB_out <=  "00011101";
    when "01111000" => SB_out <=  "10111100";
    when "10011001" => SB_out <=  "11101110";
    when "01000011" => SB_out <=  "00011010";
    when "11010110" => SB_out <=  "11110110";
    when "00001010" => SB_out <=  "01100111";
    when "00110011" => SB_out <=  "11000011";
    when "01100100" => SB_out <=  "01000011";
    when "00100001" => SB_out <=  "11111101";
    when others => SB_out <=  "00000000"; 
    end case;
  end process;
end Behavioral;
